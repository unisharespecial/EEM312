TITLE R1=1K f=1K

.model D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p 
+ M=.55 VJ=.75 FC=.5 BV=100 IBV=100u TT=11.07n)

VIN 1 0 PULSE(-10 10 0 0 0 50us 0.1ms)
VDC 3 0 DC 5

R1  1 2 1K

D2  3 2 D1N4148

D1  0 2 D1N4148

C  2 0 5nf

.control 

tran 10ns 0.5ms
plot V(1) V(2) 

.endc
.end