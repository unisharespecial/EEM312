*Soru 2 a

.MODEL MOSN NMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0
+ UO = 650 ETA = 3.0E-6 THETA = 0.1
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3
+ RSH = 0 NFS = 1E12 TPG = 1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

M1 3 1 0 2 MOSN W=90u L=1u NRS=0.333 NRD=0.333
+ AD=6.5p PD=9.0u AS=6.5p PS=9.0u

VIN 1 0 0V pulse(0V 5V 0 1ns 1ns 50ns 100ns)
VDD 3 0 5V
VBS 2 0 0V

.control
dc VDD 0V 2V 0.1V VIN 0.2V 2V 0.2V
plot -VDD#branch vs v(3)
.endc