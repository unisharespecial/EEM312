erdem

.MODEL MOSN NMOS LEVEL=2 LD=0.15U TOX=200.0E-10 
+ NSUB=5.36726E+15 VTO=0.743469 KP=8.00059E-05 GAMMA=0.543 
+ PHI=0.6 U0=655.881 UEXP=0.157282 UCRIT=31443.8 
+ DELTA=2.39824 VMAX=55260.9 XJ=0.25U LAMBDA=0.0367072 
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=1.0 RSH=70.00 
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0003 MJ=0.6585 
+ CJSW=8.0E-10 MJSW=0.2402 PB=0.58 

.MODEL MOSP PMOS LEVEL=2 LD=0.15U TOX=200.0E-10 
+ NSUB=4.3318E+15 VTO=-0.738861 KP=2.70E-05 GAMMA=0.58 
+ PHI=0.6 U0=261.977 UEXP=0.323932 UCRIT=65719.8 
+ DELTA=1.79192 VMAX=25694 XJ=0.25U LAMBDA=0.0612279 
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=-1.0 RSH=120.6 
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0005 MJ=0.5052 
+ CJSW=1.349E-10 MJSW=0.2417 PB=0.64

.subckt ters 1 2 3
M2 2 1 3 3 MOSP W=5.4u L=1.2u

M1 2 1 0 0 MOSN W=1.8u L=1.2u
.ends

Vs 3 0 3.2
Xters1 1 2 3 ters
C1 2 0 100f
Xters2 2 4 3 ters
C2 4 0 100f
Xters3 4 5 3 ters
C3 5 0 100f
Xters4 5 6 3 ters
C4 6 0 100f
Xters5 6 1 3 ters
C5 1 0 100f

.control
tran 0.1ns 60ns 0.01ns
plot v(2)
plot v(4)
plot v(5)
plot v(6)
plot v(1)
.endc
.end