**
.MODEL PMOS PMOS LEVEL = 3 
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.6
+ PHI = 0.7 VTO = -0.9 DELTA = 0.1 
+ UO = 250 ETA = 0 THETA = 0.1 
+ KP = 40E-6 VMAX = 5E4 KAPPA = 1 
+ RSH = 0 NFS = 1E12 TPG = -1 
+ XJ = 500E-9 LD = 100E-9 
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10 
+ CJ = 400E-6 PB = 1 MJ = 0.5 
+ CJSW = 300E-12 MJSW = 0.5

M2 4 1 2 3 PMOS W=1.8u L=1.2u NRS=0.333 NRD=0.333 
+ AD=6.5p PD=9.0u AS=6.5p PS=9.0u 
VIN 0 1 2
Vdd 0 2 5
Vbs 0 3 0
Vsamp 4 0 0
.control
Alter M2 W=1.8u
dc Vdd 0 5 0.1
let c1=vsamp#branch
Alter M2 W=3.6u
dc Vdd 0 5 0.1
let c2=vsamp#branch
Alter M2 W=7.2u
dc Vdd 0 5 0.1
let c3=vsamp#branch
dc Vdd 0 5 0.1
plot c1 vs v(2) c2 vs v(2) c3 vs v(2)
.endc
