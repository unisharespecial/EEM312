*20393031 Y2 soru 4 R1=1K f=1K

.model D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p 
+ M=.55 VJ=.75 FC=.5 BV=100 IBV=100u TT=11.07n)

VIN 1 0 PULSE(-10 10 0NS 2NS 2NS 0.05ms 0.1ms)
VDC 3 0 DC 5
R1  1 2 1K
D2  2 3 D1N4148
D1  2 0 D1N4148
CL  2 0 5nf

.control 

tran 20ns 0.5ms
plot V(2) 

.endc
