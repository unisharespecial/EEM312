*20294004 4. soru R1=1K f=1K

.model D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p 
+ M=.55 VJ=.75 FC=.5 BV=100 IBV=100u TT=11.07n)
VIN 1 0 PULSE(-10 10 0NS 0NS 0NS 50us 100us)
VDC 3 0 DC 5
R1  1 2 1K
D2  2 3 D1N4148
D1  0 2 D1N4148
CL  2 0 5nf
.control 
tran 10ns 500us
plot  v(1) V(2) 
.endc
