*deniz xor gate

.MODEL MOSN NMOS LEVEL=2 LD=0.15U TOX=200.0E-10 
+ NSUB=5.36726E+15 VTO=0.743469 KP=8.00059E-05 GAMMA=0.543 
+ PHI=0.6 U0=655.881 UEXP=0.157282 UCRIT=31443.8 
+ DELTA=2.39824 VMAX=55260.9 XJ=0.25U LAMBDA=0.0367072 
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=1.0 RSH=70.00 
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0003 MJ=0.6585 
+ CJSW=8.0E-10 MJSW=0.2402 PB=0.58 

.MODEL MOSP PMOS LEVEL=2 LD=0.15U TOX=200.0E-10 
+ NSUB=4.3318E+15 VTO=-0.738861 KP=2.70E-05 GAMMA=0.58 
+ PHI=0.6 U0=261.977 UEXP=0.323932 UCRIT=65719.8 
+ DELTA=1.79192 VMAX=25694 XJ=0.25U LAMBDA=0.0612279 
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=-1.0 RSH=120.6 
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0005 MJ=0.5052 
+ CJSW=1.349E-10 MJSW=0.2417 PB=0.64

M1 5 1 4 4 MOSP W=5.4u L=1.2u

M2 3 2 1 4 MOSP W=5.4u L=1.2u

M3 3 1 2 4 MOSP W=5.4u L=1.2u

M4 5 1 0 0 MOSN W=1.8u L=1.2u

M5 2 5 3 0 MOSN W=1.8u L=1.2u

M6 3 2 5 0 MOSN W=1.8u L=1.2u
vdd 4 0 5V
Vin 1 0 pulse(0V 5V 0 0ns 0ns 100ns 200ns)
Vin1 2 0 pulse(0V 5V 0 0ns 0ns 200ns 400ns)

.control
tran 0.05n 400n
plot v(3)
plot v(1)
plot v(2)
 
.endc
.end
