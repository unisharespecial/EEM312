*dcolak

.MODEL NMOSFET NMOS(VTO=1 KP=20U GAMMA=0.37 PHI=0.6 CBD=3.1E-15  CBs=3.1E-15)
M1 2 1 0 0 NMOSFET L=5U W=10U
R1 3 2 50K
C1 2 0 1P
VDC 3 0 DC 3
VIN 1 0 PULSE(0 5 0NS 2NS 2NS 500NS 1US)
.control

dc VIN 0 5 0.1

plot V(2) vs V(1)
   .endc
   .end
