*20393031 Y2 Reverse Recovery time R1=1K f=100K

.model D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p 
+ M=.55 VJ=.75 FC=.5 BV=100 IBV=100u TT=11.07n)

VIN 1 0 PULSE(0 5 0NS 2NS 2NS 0.005ms 0.01ms)
D1 1 2 D1N4148
R1 2 0 1k

.control 

tran 20ns 0.1ms
plot V(2) 

.endc
