*engin

.MODEL MOSN NMOS LEVEL = 3 
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5 
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0 
+ UO = 650 ETA = 3.0E-6 THETA = 0.1 
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3 
+ RSH = 0 NFS = 1E12 TPG = 1 
+ XJ = 500E-9 LD = 100E-9 
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10 
+ CJ = 400E-6 PB = 1 MJ = 0.5 
+ CJSW = 300E-12 MJSW = 0.5

M1 1 2 3 4 MOSN W=90u L=1u NRS=0.333 NRD=0.333 
+ AD=6.5p PD=9.0u AS=6.5p PS=9.0u

vin 2 0 0v
vdd 5 0 0v
vss 3 0 0v
vbs 4 3 0v
vsam 5 1 0v

.control

dc vdd 0 2 0.1 vin 0.2 2 0.1
plot vsam#branch vs v(1)

.endc
.end