*umut

VDC 3 0 DC 5
VIN 1 0 PULSE(0 5 0 2NS 2NS 504NS 1US)
C1 2 0 1PF
R1 3 2 50K
M1 2 1 0 0 M1 L=5U W=10U
.MODEL M1 NMOS (VTO=1 KP=20U GAMMA=0.37 PHI=0.6  CBD=3.1E-15 CBS=3.1E-15)
.DC VIN 0 5 0.01
.TRAN 0.1NS 1US
.PLOT DC V(2) VS V(1)
.PLOT TRAN V(2) V(1)
.END