netlist

VDC 3 0 DC 5
VIN 1 0 PULSE(0 5 0 2NS 500NS 1US)
R1 3 2 50K
C1 2 0 1PF
M1 2 1 0 0 M1 L=5U W=10U

.MODEL M1 NMOS(VTO=1 KP=20U GAMMA=0.37 PHI=0.6 + CBD=3.1E-15 CBS=3.1E-15)

.DC VIN 0 5 0.01
.TRAN 0.1NS 1US

.PLOT DC v(2) VS V(1)
.PLOT TRAN V(2) V(1)

.END