**

.MODEL D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p + M=.55 VJ=.75 FC=.5 BV=50 IBV= 100u TT=11.07n)
D1 1 2 D1N4148
R1 2 0 10K
Vin 1 0 5V DC
.control

DC Vin -300 200 0.1
plot -Vin#branch vs v(1)-v(2)
.endc
.end
