**

.MODEL D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p + M=.55 VJ=.75 FC=.5 BV=100 IBV= 100u TT=11.07n)
D1 2 0 D1N4148
D2 2 3 D1N4148
R1 1 2 1K
C 2 0 5nf
Vin 1 0 PULSE (-10 10 0NS 2NS 2NS 0.05ms 0.1ms)
VDD 3 0 5V

.control
tran 1ns 0.5ms
plot V(2) 
.endc
.end
