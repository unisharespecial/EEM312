*Soru 4

VDD 3 0 DC 5
VIN 1 0 PULSE(-10 10 0 0 0 50us 100us)
R1  1 2 1K
D1  2 3 D1N4148
D2  0 2 D1N4148
C   2 0 5NF

	
.model D1N4148 D(IS=5.84n N=1.94 RS=.7017 XTI=3 EG=1.11 CJO=.95p 
+ M=.55 VJ=.75 FC=.5 BV=100 IBV=100u TT=11.07n)


.CONTROL

TRAN 10ns 500us

PLOT V(1)  V(2)
.ENDC 


.END
     