* Ugur Zongur 20395080
* Lab: Software #5

.MODEL MOSN NMOS LEVEL=2 LD=0.15U TOX=200.0E-10
+ NSUB=5.36726E+15 VTO=0.743469 KP=8.00059E-05 GAMMA=0.543
+ PHI=0.6 U0=655.881 UEXP=0.157282 UCRIT=31443.8
+ DELTA=2.39824 VMAX=55260.9 XJ=0.25U LAMBDA=0.0367072
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=1.0 RSH=70.00
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0003 MJ=0.6585
+ CJSW=8.0E-10 MJSW=0.2402 PB=0.58

.MODEL MOSP PMOS LEVEL=2 LD=0.15U TOX=200.0E-10
+ NSUB=4.3318E+15 VTO=-0.738861 KP=2.70E-05 GAMMA=0.58
+ PHI=0.6 U0=261.977 UEXP=0.323932 UCRIT=65719.8
+ DELTA=1.79192 VMAX=25694 XJ=0.25U LAMBDA=0.0612279
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=-1.0 RSH=120.6
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0005 MJ=0.5052
+ CJSW=1.349E-10 MJSW=0.2417 PB=0.64

M1 3 1 0 0 MOSN W=19.66um L=1um NRS=0.323 NRD=0.323
+ AD=15p PD=17.4u AS=15p PS=17.5u

M2 3 1 2 2 MOSP W=57.8u L=1um NRS=0.129 NRD=0.129
+ AD=38.75p PD=36u AS=38.75p PS=36u

CL 3 0 1pF

* V1=0, V2=3.2V, td=0, tr=tf=1n, pw=50n, per=100n
VIN 1 0 0V pulse(0V 3.2V 0 1ns 1ns 50ns 100ns)
VDD 2 0 3.2V

.control

* dc VIN 0 3.2 0.1
* plot v(3) vs v(1) v(1) vs v(1)


tran 0.1ns 100ns
plot v(3) v(1)

.endc