s1


.MODEL MOSN NMOS LEVEL=2 LD=0.15U TOX=200.0E-10 
+ NSUB=5.36726E+15 VTO=0.743469 KP=8.00059E-05 GAMMA=0.543 
+ PHI=0.6 U0=655.881 UEXP=0.157282 UCRIT=31443.8 
+ DELTA=2.39824 VMAX=55260.9 XJ=0.25U LAMBDA=0.0367072 
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=1.0 RSH=70.00 
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0003 MJ=0.6585 
+ CJSW=8.0E-10 MJSW=0.2402 PB=0.58 

.MODEL MOSP PMOS LEVEL=2 LD=0.15U TOX=200.0E-10 
+ NSUB=4.3318E+15 VTO=-0.738861 KP=2.70E-05 GAMMA=0.58 
+ PHI=0.6 U0=261.977 UEXP=0.323932 UCRIT=65719.8 
+ DELTA=1.79192 VMAX=25694 XJ=0.25U LAMBDA=0.0612279 
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=-1.0 RSH=120.6 
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0005 MJ=0.5052 
+ CJSW=1.349E-10 MJSW=0.2417 PB=0.64

*  D G S B

M1 3 2 1 1 MOSP W=3.6u L=1.2u
M2 2 4 5 5 MOSP W=3.6u L=1.2u
M3 4 2 5 5 MOSP W=3.6u L=1.2u

M4 3 2 0 0 MOSN W=1.8u L=1.2u
M5 3 4 5 5 MOSN W=1.8u L=1.2u
M6 5 3 4 4 MOSN W=1.8u L=1.2u

vdd 1 0 5V
v2 2 0 0v
v4 4 0 0v

*Vin1 2 0 pulse(0V 5V 0 0ns 0ns 100ns 200ns)
*Vin2 4 0 pulse(0V 5V 0 0ns 0ns 200ns 400ns)

.control
tran 0.05n 500n
plot v(2) v(4) v(5)
 
.endc
.end
