*can
.MODEL NMOS NMOS
+LEVEL = 49
+LINT = 4.E-08 TOX = 4.E-09 VTH0 = 0.3999 RDSW = 250
+LMIN=1.8E-7 LMAX=1.8E-7 WMIN=1.8E-7 WMAX=1.0E-4 TREF=27.0 VERSION =3.1
+XJ= 6.0000000E-08 NCH= 5.9500000E+17
+LLN= 1.0000000 LWN= 1.0000000 WLN= 0.00 WWN= 0.00 LL= 0.00
+LW= 0.00 LWL= 0.00 WINT= 0.00 WL= 0.00 WW= 0.00 WWL= 0.00
+MOBMOD= 1 BINUNIT= 2 XL= 0
+XW= 0 BINFLAG= 0 DWG= 0.00 DWB= 0.00
+K1= 0.5613000 K2= 1.0000000E-02
+K3= 0.00 DVT0= 8.0000000 DVT1= 0.7500000
+DVT2= 8.0000000E-03 DVT0W= 0.00 DVT1W= 0.00
+DVT2W= 0.00 NLX= 1.6500000E-07 W0= 0.00
+K3B= 0.00 NGATE= 5.0000000E+20
+VSAT= 1.3800000E+05 UA= -7.0000000E-10 UB= 3.5000000E-18
+UC= -5.2500000E-11 PRWB= 0.00
+PRWG= 0.00 WR= 1.0000000 U0= 3.5000000E-02
+A0= 1.1000000 KETA= 4.0000000E-02 A1= 0.00
+A2= 1.0000000 AGS= -1.0000000E-02 B0= 0.00 B1= 0.00
+VOFF= -0.12350000 NFACTOR= 0.9000000 CIT= 0.00
+CDSC= 0.00 CDSCB= 0.00 CDSCD= 0.00
+ETA0= 0.2200000 ETAB= 0.00 DSUB= 0.8000000
+PCLM= 5.0000000E-02 PDIBLC1= 1.2000000E-02 PDIBLC2= 7.5000000E-03
+PDIBLCB= -1.3500000E-02 DROUT= 1.7999999E-02 PSCBE1= 8.6600000E+08
+PSCBE2= 1.0000000E-20 PVAG= -0.2800000 DELTA= 1.0000000E-02
+ALPHA0= 0.00 BETA0= 30.0000000
+KT1= -0.3700000 KT2= -4.0000000E-02 AT= 5.5000000E+04
+UTE= -1.4800000 UA1= 9.5829000E-10 UB1= -3.3473000E-19
+UC1= 0.00 KT1L= 4.0000000E-09 PRT= 0.00
+CJ= 0.00365 MJ= 0.54 PB= 0.982
+CJSW= 7.9E-10 MJSW= 0.31 PHP= 0.841
+CTA= 0 CTP= 0 PTA= 0
+PTP= 0 JS=1.50E-08 JSW=2.50E-13
+N=1.0 XTI=3.0 CGDO=2.786E-10
+CGSO=2.786E-10 CGBO=0.0E+00 CAPMOD= 2
+NQSMOD= 0 ELM= 5 XPART= 1
+CGSL= 1.6E-10 CGDL= 1.6E-10 CKAPPA= 2.886
+CF= 1.069E-10 CLC= 0.0000001 CLE= 0.6
+DLC= 4E-08 DWC= 0 VFBCV= -1
M1 3 1 0 2 NMOS W=5u L=0.18u NRS=0.333 NRD=0.333
+ AD=6.5p PD=9.0u AS=6.5p PS=9.0u
VIN 1 0 1
VDD 3 0 5
VBS 2 0 0
.control
dc VDD 0 2 0.1 VIN 0.2 2 0.2 
plot -VDD#branch vs v(3)
.endc
