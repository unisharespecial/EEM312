*
R1 1 2 50K
C1 2 0 1P
VIN 3 0 PULSE(0 5 0 2NS 2NS 504NS 1US)
VDC 1 0 DC 3
.MODEL NMOSFET NMOS(VTO=1 KP=20U GAMMA=0.37 PHI=0.6  CBD=3.1E-15  CBS=3.1E-15)
M1 2 3 0 0 NMOSFET L=5U W=10U
*.DC VIN 0 10 0.1
.TRAN 0.1nS 2US
*.PLOT DC v(2)
.PLOT TRAN V(2) V(3)
.END