*NMOS TERSLEYICI
R1 1 2 100K
C1 2 0 1ff
VIN 3 0 PULSE(0 5 0NS 2NS 2NS 500NS 1US)
VDC 1 0 DC 3.1

.MODEL MOSN NMOS LEVEL=2 LD=0.15U TOX=200.0E-10
+ NSUB=5.36726E+15 VTO=0.743469 KP=8.00059E-05 GAMMA=0.543
+ PHI=0.6 U0=655.881 UEXP=0.157282 UCRIT=31443.8
+ DELTA=2.39824 VMAX=55260.9 XJ=0.25U LAMBDA=0.0367072
+ NFS=1E+12 NEFF=1.001 NSS=1E+11 TPG=1.0 RSH=70.00
+ CGDO=4.3E-10 CGSO=4.3E-10 CJ=0.0003 MJ=0.6585
+ CJSW=8.0E-10 MJSW=0.2402 PB=0.58

M1 2 3 0 0 MOSN W=1.8U L=1.2U NRS=0.333 NRD=0.333
+ AD=6.5P PD=9.0U AS=6.5P PS=9.0U



.CONTROL

DC VIN 0 5 0.1 
PLOT V(2) VS V(3)

.ENDC