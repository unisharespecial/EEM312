BSIM3V3 MODEL�

.model MOSN NMOS
+Level= 8
+Tnom=27.0 Nch= 2.498E+17 Tox=9E-09 Xj=1.00000E-07
+Lint=9.36e-8 Wint=1.47e-7 Vth0= .6322 K1= .756 K2= -3.83e-2 K3= -2.612
+Dvt0= 2.812 Dvt1= 0.462 Dvt2=-9.17e-2
+Nlx= 3.52291E-08 W0= 1.163e-6 K3b= 2.233
+Vsat= 86301.58 Ua= 6.47e-9 Ub= 4.23e-18 Uc=-4.706281E-11
+Rdsw= 650 U0= 388.3203 wr=1 A0= .3496967 Ags=.1 B0=0.546 B1= 1
+ Dwg = -6.0E-09 Dwb = -3.56E-09 Prwb = -.213
+Keta=-3.605872E-02 A1= 2.778747E-02 A2= .9
+Voff=-6.735529E-02 NFactor= 1.139926 Cit= 1.622527E-04
+Cdsc=-2.147181E-05 Cdscb= 0 Dvt0w = 0 Dvt1w = 0 Dvt2w = 0
+ Cdscd = 0 Prwg = 0 Eta0= 1.0281729E-02 Etab=-5.042203E-03
+Dsub= .31871233 Pclm= 1.114846 Pdiblc1= 2.45357E-03 Pdiblc2= 6.406289E-03
+Drout= .31871233 Pscbe1= 5000000 Pscbe2= 5E-09 Pdiblcb = -.234
+Pvag= 0 delta=0.01 Wl = 0 Ww = -1.420242E-09 Wwl = 0
+ Wln = 0 Wwn = .2613948 Ll = 1.300902E-10
+ Lw = 0 Lwl = 0 Lln = .316394 Lwn = 0 kt1=-.3 kt2=-.051
+At= 22400 Ute=-1.48
+Ua1= 3.31E-10 Ub1= 2.61E-19 Uc1= -3.42e-10 Kt1l=0 Prt=764.3

M1 2 1 3 5 MOSN W=10u L=2u NRS=0.333 NRD=0.333
+ AD=6.5p PD=9.0u AS=6.5p PS=9.0u

R1 2 4 10k
Vsamp  3 0 0
Vdd  4 0 5
VIN  1 0 5
Vbs 5 0 0

.control

dc Vdd 0 3 0.1 VIN 0 3 0.1
plot Vsamp#branch vs V(2)

.endc
.end




